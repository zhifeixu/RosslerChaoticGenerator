library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


package nn_package is

    -- Network architecture parameters
    constant NUM_X : integer := 3; -- Number of inputs
    constant NUM_L1 : integer := 20; -- Number of hidden layer neurons
    constant NUM_Y : integer := 3; -- Number of outputs
    
    -- Data representation constants
    constant N : integer := 32; -- Number of bits (data width)
    constant F : integer := 14; -- Number of fractional bits
    constant I : integer := N-F; -- Number of integer bits
    constant ONE : real := 2.0**F;
    constant ONE_int : integer := integer(ONE); -- 1 in fixed point representation
    
    -- Array types (for representing signals throughout the network
    type x_array is array(0 to NUM_X-1) of signed(N-1 downto 0); -- Array of inputs
    type y_array is array(0 to NUM_Y-1) of signed(N-1 downto 0); -- Array of outputs
    type sum1_array is array(0 to NUM_L1-1) of signed(N-1 downto 0); -- Array of hidden neuron outputs
    type sum2_array is array(0 to NUM_Y-1) of signed(N-1 downto 0); -- Array of output neuron outputs
    type a_array is array(0 to NUM_L1-1) of signed(N-1 downto 0); -- Array of hidden activation function outputs
    
    -- Array types (real valued for representation of bias, weight and
    -- normalization parameters
    type b1r_array is array(0 to NUM_L1-1) of real; -- Hidden layer biases
    type b2r_array is array(0 to NUM_Y-1) of real; -- Output layer biases
    type w1r_array is array(0 to NUM_X*NUM_L1-1) of real; -- Hidden layer weights
    type w2r_array is array(0 to NUM_L1*NUM_Y-1) of real; -- Output layer weights
    type p1r_array is array(0 to NUM_X-1) of real; -- Normalization parameters
    type p2r_array is array(0 to NUM_Y-1) of real; -- Denormalization parameters

    -- Array types (signed valued for representation of bias, weight and
    -- normalization parameters
    type b1_array is array (0 to NUM_L1-1) of signed(N-1 downto 0); -- Hidden layer biases
    type b2_array is array (0 to NUM_Y-1) of signed(N-1 downto 0); -- Output layer biases
    type w1_array is array (0 to NUM_L1-1) of x_array; -- Hidden layer weights
    type w2_array is array (0 to NUM_Y-1) of a_array; -- Output layer weights
    type p1_array is array (0 to NUM_X-1) of signed(N-1 downto 0); -- Normalization parameters
    type p2_array is array (0 to NUM_Y-1) of signed(N-1 downto 0); -- Denormalization parameters
    
    -- Real weights and biases
    -- hidden layer biases
    constant b1r : b1r_array := (4.1017041891290695332,-3.509108718728506382,3.3246597636241888019,-2.1699268616627671591,3.2542397371625528812,-1.5093288425161139887,0.62634630231450028059,1.4732014703897955421,0.27094695152384584702,-0.10258621270142366522,0.026875628244393112015,1.1046732460802590747,0.15962048163824224534,1.6242783487012899535,1.7790059428500684113,3.4916440834872006782,1.4356841189530271663,-4.3697872061953484391,-4.3821388062575792333,2.9681886535512580494); 
    -- output layer biases
    constant b2r : b2r_array := (-0.59281491019938892251,-0.051035225522110011509,-0.32588867388349657128); 
    -- hidden layer weights
    constant w1r : w1r_array := (-1.2052508491243405508,2.5350766791781320642,-2.3001454218868060408,1.5028882343963589907,-2.1680779705668995483,2.3759234047540878088,-1.2689167957106335383,2.4261332335130552096,-2.3246474765384190775,1.6683563383562514115,-2.5919038144030288606,-0.59038287913994025313,-3.0304320573760787916,-0.87103255122977474301,-1.1675438895168368525,1.0946126898434294095,-2.0537419686507352168,1.2702965112400921299,-0.27631269028288085732,-0.016625060996039872641,-0.32247457266110646223,-0.49034081230074116897,-0.030114091344010981977,0.60286466339608979492,-1.2881797525505771507,-1.1073583162560693971,3.1255556111717446299,0.10901064764612625191,0.1417255234788266649,0.064672621860391327209,0.35506651064334399104,0.025707398588206777784,-0.43360434145735987643,1.4956306310369502643,1.0097288083786926105,-3.1029395290484087511,0.11299252645790139327,-0.2146327564620602868,0.16726776733802981023,2.0759977986302291519,0.5776694041639371946,-2.3754520021797405072,2.2612467525587187644,0.72469423107150610086,-2.6082824730286593429,1.7600817673256878848,1.323112593297646411,-2.2936992564295648478,0.47622144013422268438,0.64553591937648946431,0.21581513923212128359,-0.51909382575176732377,2.3504537011129560398,1.801089403491407559,-1.3123511607542879265,2.2197649661470921778,2.2069273035839311881,0.69693542153956244967,-1.3484867539374156831,1.0112396847431439628); 
    -- output layer weights
    constant w2r : w2r_array := (-0.47921955871658555859,0.37331482257153880688,0.60318174400441981753,0.0011696899793432983129,-0.013013155234985128786,0.020312715811731250209,0.023356094187708818094,-0.5632857952630990761,0.00096572720395745627591,2.8225719532555197944,1.0795641210511286445,-0.0047958183787715985905,2.0969290315422237647,0.29827614443142014267,-0.33129982747158925882,0.79481986701836770948,0.08245384736040037299,0.32752052381503848899,-0.7525349329287929212,0.02720385068496215808,-0.13634835555153831943,-0.24311412136193039091,-0.3349077731797108215,-0.0014058527909256099148,0.016905672663166976255,-0.020893570461050000459,-0.016275771962094839201,0.15225921061572333937,0.00016153157055105813594,3.6118161306903107111,-0.28269261161968056717,0.0031623152116082653765,-2.2726527284609816526,-0.0071649349189385688752,-0.018018785332376729275,0.68984106633904362926,0.11562997347958314798,-0.23616097273072594875,0.12098761090038097354,-0.03061851962328921567,0.26264162355182169017,0.13211993295477106325,0.081174896988630937389,0.00061121955348588069383,-0.017624204700736511436,0.0075848837229339511473,-1.4103180448264980296,0.79259308702159925186,-0.0021388125994798528294,1.2602387325624233583,-0.71094508689594548834,0.0021066777542095862195,0.76437005547281478002,0.069970791467323753543,-0.091725944007985532602,-0.21528980965343263998,0.041744117925318791062,-0.2549055702521065836,-0.082128541161245682822,0.0085879024479075215248); 
    
    -- Parameters for input and output processing
    -- min inputs
    constant p11r : p1r_array := (0.0, 0.0, 0.0); 
    -- 2/(max inputs - min inputs)
    constant p12r : p1r_array := (2.0,2.0,2.0); -- 2/(max - min) = 2/(1 - 0) == 2
    -- 1's array
    constant p13r : p1r_array := (1.0000000000, 1.0000000000, 1.0000000000); 
    
    -- 1's array
    constant p21r : p2r_array := (1.0000000000, 1.0000000000, 1.0000000000);
    -- (max targets - min targets)/2
    constant p22r : p2r_array := (0.5, 0.5, 0.5); -- = (1-0)/2 == 0.5
    -- min targets
    constant p23r : p2r_array := (0.0, 0.0, 0.0);

end package nn_package;

